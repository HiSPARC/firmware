-- EASE/HDL begin --------------------------------------------------------------
-- Architecture 'a0' of 'DUMMIES.
--------------------------------------------------------------------------------
-- Copy of the interface declaration of Entity 'DUMMIES' :
-- 
--   port(
--     ADC_1_NEG_OR : in     std_logic;
--     ADC_1_POS_OR : in     std_logic;
--     ADC_2_NEG_OR : in     std_logic;
--     ADC_2_POS_OR : in     std_logic;
--     LED4         : out    std_logic;
--     LED5         : out    std_logic;
--     LED6         : out    std_logic;
--     LED7         : out    std_logic;
--     LED8         : out    std_logic;
--     LED9         : out    std_logic);
-- 
-- EASE/HDL end ----------------------------------------------------------------

architecture a0 of DUMMIES is

begin

-- The ADC input signals are not connected

-- LED1 is used for SLAVE_PRESENT
-- LED2 is used for MASTER (GPS PRESENT)
-- LED3 is used for COINC
  LED4 <= '1';
  LED5 <= '1';
  LED6 <= '1';
  LED7 <= '1';
  LED8 <= '1';
  LED9 <= '1';

end architecture a0 ; -- of DUMMIES

